module control_state(

);

//boilerplate