module control_unit(

);

//boilerplate for sequential control unit

//top level -> control state + control logic 