module program_counter(

);

//boilerplate