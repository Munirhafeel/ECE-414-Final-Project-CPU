module instruction_register(

);

//boiler plate for IR